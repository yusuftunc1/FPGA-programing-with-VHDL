library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

